module _nand(input a, input b, output c);
assign c = ~(a & b);
endmodule

